netcdf SAR_drift_data {
dimensions:
    time = UNLIMITED ;
    x = 361 ;
    y = 361 ;

variables: 
    float Speed_kmdy(time, y, x) ;
        Speed_kmdy:long_name = "Speed in km/day" ;
		Speed_kmdy:standard_name = "sea_ice_speed" ;
        Speed_kmdy:ioos_category = "SAR daily sea-ice drift" ;
        Speed_kmdy:units = "km/day" ;
        Speed_kmdy:grid_mapping = "spatial_ref" ;


    float U_vel_ms(time, y, x) ;
        U_vel_ms:long_name = "Zonal Velocity" ;
		U_vel_ms:standard_name = "movement_in_x_direction" ;
        U_vel_ms:ioos_category = "SAR daily sea-ice drift" ;
        U_vel_ms:units = "m/s" ;
        U_vel_ms:grid_mapping = "spatial_ref" ;


    float V_vel_ms(time, y, x) ;
        V_vel_ms:long_name = "Meridional Velocity" ;
		V_vel_ms:standard_name = "movement_in_y_direction" ;		
        V_vel_ms:ioos_category = "SAR daily sea-ice drift" ;
        V_vel_ms:units = "m/s" ;
        V_vel_ms:grid_mapping = "spatial_ref" ;


    float Bear_deg(time, y, x) ;
        Bear_deg:long_name = "Bearing" ;
		Bear_deg:standard_name = "direction_true_north" ;
        Bear_deg:ioos_category = "SAR daily sea-ice drift" ;
        Bear_deg:units = "degrees" ;
        Bear_deg:grid_mapping = "spatial_ref" ;


    float x(x) ;
        x:actual_range = 0.0, 0.0;
        x:axis = "X" ;
        x:comment = "x values are the centers of the grid cells" ;
        x:ioos_category = "Location" ;
        x:long_name = "x coordinate of projection" ;
        x:standard_name = "projection_x_coordinate" ;
        x:units = "m" ;

    float y(y) ;
        y:actual_range = 0.0, 0.0 ;
        y:axis = "Y" ;
        y:comment = "y values are the centers of the grid cells" ;
        y:ioos_category = "Location" ;
        y:long_name = "y coordinate of projection" ;
        y:standard_name = "projection_y_coordinate" ;
        y:units = "m" ;

    double time(time) ;
        time:actual_range = 1712793600.0, 1712880000.0 ;
        time:axis = "T" ;
        time:comment = "This is the 00Z reference time. Note that products are nowcasted to be valid specifically at the time given here." ;
        time:CoordinateAxisType = "Time" ;
        time:ioos_category = "Time" ;
        time:long_name = "Centered Time" ;
        time:standard_name = "time" ;
        time:time_origin = "01-Jan-1970 0:00:00" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;


// global attributes:
	:acknowledgement = "Produced by NOAA using IABP data." ;
	:cdm_data_type = "Grid" ;
	:contributor_name = "NOAA PolarWatch, Southwest Fisheries Science Center, NESDIS STAR, U.S. National Ice Center" ;
	:contributor_role = "Producer, Publisher, Advisor, Originator" ;
	:Conventions = "CF-1.8, ACDD-1.3" ;
	:creator_email = "brendon.gory@noaa.gov" ;
	:creator_institution = "CIRA/NOAA" ;
	:creator_name = "Brendon Gory" ;
	:creator_type = "Institution" ;
	:creator_url = "https://noaa.gov/" ;
	:date_created = "FILL_DATE_CREATED" ;
	:grid_mapping__ChunkSizes = 1 ;
	:grid_mapping_false_easting = 0 ;
	:grid_mapping_false_northing = 0 ;
	:grid_mapping_latitude_of_projection_origin = 90 ;
	:grid_mapping_name = "polar_stereographic" ;
	:grid_mapping_proj4text = "+proj=stere +lat_0=90 +lat_ts=60 +lon_0=-80 +k=1 +x_0=0 +y_0=0 +a=6378137 +b=6356257 +units=m +no_defs" ;
	:grid_mapping_semi_major_axis = 6378137 ;
	:grid_mapping_semi_minor_axis = 6356257 ;
	:grid_mapping_spatial_ref = "PROJCS[\"unknown\",GEOGCS[\"unknown\",DATUM[\"unknown\",SPHEROID[\"unknown\",6378137,291.505347349177]],PRIMEM[\"Greenwich\",0,AUTHORITY[\"EPSG\",\"8901\"]],UNIT[\"degree\",0.0174532925199433,AUTHORITY[\"EPSG\",\"9122\"]]],PROJECTION[\"Polar_Stereographic\"],PARAMETER[\"latitude_of_origin\",60],PARAMETER[\"central_meridian\",-80],PARAMETER[\"false_easting\",0],PARAMETER[\"false_northing\",0],UNIT[\"metre\",1,AUTHORITY[\"EPSG\",\"9001\"]],AXIS[\"Easting\",SOUTH],AXIS[\"Northing\",SOUTH]]" ;
	:grid_mapping_standard_parallel = 60 ;
	:grid_mapping_straight_vertical_longitude_from_pole = -80 ;
	:grid_mapping_units = "m" ;
	:history = "02 Apr 2025: First version of convert SAR dailt drift to NetCDF" ;
	:infoUrl = "https://coastwatch.noaa.gov/cwn/products/sar-composite-arctic-imagery-normalized-radar-cross-section.html" ;
	:institution = "NOAA CoastWatch" ;
	:instrument = "See website for detailshttps://coastwatch.noaa.gov/cwn/products/sar-composite-arctic-imagery-normalized-radar-cross-section.html" ;
	:keywords = "Earth Science > Cryosphere > Sea Ice > Ice Extent, Earth Science > Cryosphere > Snow/Ice > Snow Cover, GEOGRAPHIC REGION > ARCTIC, GEOGRAPHIC REGION > NORTHERN HEMISPHERE, GEOGRAPHIC REGION > POLAR" ;
	:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Keywords, Version 9.0" ;
	:license = "U.S. Government Work (public domain)" ;
	:metadata_link = "https://coastwatch.noaa.gov/cwn/products/sar-composite-arctic-imagery-normalized-radar-cross-section.html" ;
	:naming_authority = "gov.noaa.polarwatch" ;
	:ncei_template_version = "NCEI_NetCDF_Grid_Template_v2.0" ;
	:platform = "Earth Observation Satellites, In Situ Land-based Platforms, Ground Stations, Models/Analyses" ;
	:platform_vocabulary = "NASA Global Change Master Directory (GCMD) Keywords, Version 9.0" ;
	:processing_level = "NOAA Level 4" ;
	:product_version = "Version 1" ;
	:project = "NOAA Polarwatch" ;
	:publisher_email = "coastwatch at noaa dot gov" ;
	:publisher_institution = "NOAA CoastWatch" ;
	:publisher_name = "NOAA CoastWatch" ;
	:publisher_type = "Institutional" ;
	:publisher_url = "coastwatch.noaa.gov" ;
	:references = "See website for detailshttps://coastwatch.noaa.gov/cwn/products/sar-composite-arctic-imagery-normalized-radar-cross-section.html" ;
	:source = "SAR Daily Drift dataset" ;
	:sourceUrl = "https://www.star.nesdis.noaa.gov/socd/mecb/sar/AKDEMO_products/COMPOSITE_TIFF/DRIFT_SHAPEFILES/" ;
	:standard_name_vocabulary = "CF Standard Name Table (Version 72, 10 March 2020)" ;
	:summary = "NetCDF version of the SAR Daily Drift dataset. This dataset includes the starting and ending coordinates (latitude and longitude), start and end observation dates, total distance traveled, and drift bearing over the observation period." ;
	:title = "SAR drift data converted from raw text form to NetCDF" ;
	:time_coverage_duration = "P1D" ;
	:time_coverage_resolution = "P1D" ;
	:time_coverage_end = "FILL_MAX_TIME" ;
	:time_coverage_start = "FILL_MIN_TIME" ;
}